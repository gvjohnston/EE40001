[aimspice]
[description]
1010
.MODEL CMOSN NMOS LEVEL=2 LD=0.250000U TOX=417.000008E-10
+ NSUB=6.108619E+14 VTO=0.825008 KP=4.919000E-05 GAMMA=0.172
+ PHI=0.6 UO=594 UEXP=6.682275E-02 UCRIT=5000
+ DELTA=5.08308 VMAX=65547.3 XJ=0.250000U LAMBDA=6.636197E-03
+ NFS=1.98E+11 NEFF=1 NSS=1.000000E+10 TPG=1.000000
+ RSH=32.740000 CGDO=3.105345E-10 CGSO=3.105345E-10 CGBO=3.848530E-10
+ CJ=9.494900E-05 MJ=0.847099 CJSW=4.410100E-10 MJSW=0.334060 PB=0.800000

.MODEL CMOSP PMOS LEVEL=2 LD=0.227236U TOX=417.000008E-10
+ NSUB=1.056124E+16 VTO=-0.937048 KP=1.731000E-05 GAMMA=0.715
+ PHI=0.6 UO=209 UEXP=0.233831 UCRIT=47509.9
+ DELTA=1.07179 VMAX=100000 XJ=0.250000U LAMBDA=4.391428E-02
+ NFS=3.27E+11 NEFF=1.001 NSS=1.000000E+10 TPG=-1.000000
+ RSH=72.960000 CGDO=2.822585E-10 CGSO=2.822585E-10 CGBO=5.292375E-10
+ CJ=3.224200E-04 MJ=0.584956 CJSW=2.979100E-10 MJSW=0.310807 PB=0.800000

M1 3 2 4 1 CMOSP L=2u W=25u AD=137.5p PD=61u AS=137.5p PS=61u 
* M1 DRAIN GATE SOURCE BULK (12 10 14 35) 

VB 1 0 DC 5V
VGD 2 3
VSD 4 3

[dc]
2
VSD
0V
-10V
-0.1V
VGD
-1V
-5V
-1V
[ana]
1 1
0
1 1
1 1 -8.23994E-018 0.0025
1
i(vsd)
[end]
